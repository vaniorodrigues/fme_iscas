/*
* @Author: Vanio Rodrigues Filho
* @Date:   2018-03-21 10:49:04
* @Last Modified by:   VanioRodrigues
* @Last Modified time: 2018-04-05 14:38:08
*/

//`include "register.v"

module SR_horizontal(
	clock, 
	reset,
	enable,
	enable_read,
	in_0,
	in_1,
	in_2,
	in_3,
	in_4,
	in_5,
	in_6,
	in_7,
	in_8,
	in_9,
	in_10,
	in_11,
	in_12,
	in_13,
	in_14,
	in_15,
	in_16,
	in_17,
	in_18,
	in_19,
	in_20,
	in_21,
	in_22,
	in_23,
	in_24,
	in_25,
	in_26,
	out_0,
	out_1,
	out_2,
	out_3,
	out_4,
	out_5,
	out_6,
	out_7,
	out_8,
	out_9,
	out_10,
	out_11,
	out_12,
	out_13,
	out_14,
	out_15
);

//--------------------------------- Parameters -----------------------------//

parameter DATAWIDTH = 8;

//--------------------------------- Input ports -----------------------------//

input clock, reset, enable, enable_read;

input signed [DATAWIDTH+7:0] in_0, in_1, in_2, in_3, in_4, in_5, in_6, in_7, in_8, in_9, in_10, in_11, in_12, in_13, in_14, in_15, in_16,in_17,in_18,in_19,in_20,in_21,in_22,in_23,in_24,in_25,in_26;

//--------------------------------- Output ports -----------------------------//

output reg signed [DATAWIDTH+7:0] out_0, out_1, out_2, out_3, out_4, out_5, out_6, out_7, out_8, out_9, out_10, out_11, out_12, out_13, out_14, out_15;

//--------------------------------- Internal Wires -----------------------------//

wire signed [DATAWIDTH+7:0] out_of_0_0,out_of_0_1,out_of_0_2,out_of_0_3,out_of_0_4,out_of_0_5,out_of_0_6,out_of_0_7,out_of_0_8,out_of_0_9,out_of_0_10,out_of_0_11,out_of_0_12,out_of_0_13,out_of_0_14,out_of_0_15,out_of_0_16,out_of_0_17,out_of_0_18,out_of_0_19,out_of_0_20,out_of_0_21,out_of_0_22,out_of_0_23,out_of_0_24,out_of_0_25,out_of_0_26,out_of_1_0,out_of_1_1,out_of_1_2,out_of_1_3,out_of_1_4,out_of_1_5,out_of_1_6,out_of_1_7,out_of_1_8,out_of_1_9,out_of_1_10,out_of_1_11,out_of_1_12,out_of_1_13,out_of_1_14,out_of_1_15,out_of_1_16,out_of_1_17,out_of_1_18,out_of_1_19,out_of_1_20,out_of_1_21,out_of_1_22,out_of_1_23,out_of_1_24,out_of_1_25,out_of_1_26,out_of_2_0,out_of_2_1,out_of_2_2,out_of_2_3,out_of_2_4,out_of_2_5,out_of_2_6,out_of_2_7,out_of_2_8,out_of_2_9,out_of_2_10,out_of_2_11,out_of_2_12,out_of_2_13,out_of_2_14,out_of_2_15,out_of_2_16,out_of_2_17,out_of_2_18,out_of_2_19,out_of_2_20,out_of_2_21,out_of_2_22,out_of_2_23,out_of_2_24,out_of_2_25,out_of_2_26,out_of_3_0,out_of_3_1,out_of_3_2,out_of_3_3,out_of_3_4,out_of_3_5,out_of_3_6,out_of_3_7,out_of_3_8,out_of_3_9,out_of_3_10,out_of_3_11,out_of_3_12,out_of_3_13,out_of_3_14,out_of_3_15,out_of_3_16,out_of_3_17,out_of_3_18,out_of_3_19,out_of_3_20,out_of_3_21,out_of_3_22,out_of_3_23,out_of_3_24,out_of_3_25,out_of_3_26,out_of_4_0,out_of_4_1,out_of_4_2,out_of_4_3,out_of_4_4,out_of_4_5,out_of_4_6,out_of_4_7,out_of_4_8,out_of_4_9,out_of_4_10,out_of_4_11,out_of_4_12,out_of_4_13,out_of_4_14,out_of_4_15,out_of_4_16,out_of_4_17,out_of_4_18,out_of_4_19,out_of_4_20,out_of_4_21,out_of_4_22,out_of_4_23,out_of_4_24,out_of_4_25,out_of_4_26,out_of_5_0,out_of_5_1,out_of_5_2,out_of_5_3,out_of_5_4,out_of_5_5,out_of_5_6,out_of_5_7,out_of_5_8,out_of_5_9,out_of_5_10,out_of_5_11,out_of_5_12,out_of_5_13,out_of_5_14,out_of_5_15,out_of_5_16,out_of_5_17,out_of_5_18,out_of_5_19,out_of_5_20,out_of_5_21,out_of_5_22,out_of_5_23,out_of_5_24,out_of_5_25,out_of_5_26,out_of_6_0,out_of_6_1,out_of_6_2,out_of_6_3,out_of_6_4,out_of_6_5,out_of_6_6,out_of_6_7,out_of_6_8,out_of_6_9,out_of_6_10,out_of_6_11,out_of_6_12,out_of_6_13,out_of_6_14,out_of_6_15,out_of_6_16,out_of_6_17,out_of_6_18,out_of_6_19,out_of_6_20,out_of_6_21,out_of_6_22,out_of_6_23,out_of_6_24,out_of_6_25,out_of_6_26,out_of_7_0,out_of_7_1,out_of_7_2,out_of_7_3,out_of_7_4,out_of_7_5,out_of_7_6,out_of_7_7,out_of_7_8,out_of_7_9,out_of_7_10,out_of_7_11,out_of_7_12,out_of_7_13,out_of_7_14,out_of_7_15,out_of_7_16,out_of_7_17,out_of_7_18,out_of_7_19,out_of_7_20,out_of_7_21,out_of_7_22,out_of_7_23,out_of_7_24,out_of_7_25,out_of_7_26,out_of_8_0,out_of_8_1,out_of_8_2,out_of_8_3,out_of_8_4,out_of_8_5,out_of_8_6,out_of_8_7,out_of_8_8,out_of_8_9,out_of_8_10,out_of_8_11,out_of_8_12,out_of_8_13,out_of_8_14,out_of_8_15,out_of_8_16,out_of_8_17,out_of_8_18,out_of_8_19,out_of_8_20,out_of_8_21,out_of_8_22,out_of_8_23,out_of_8_24,out_of_8_25,out_of_8_26,out_of_9_0,out_of_9_1,out_of_9_2,out_of_9_3,out_of_9_4,out_of_9_5,out_of_9_6,out_of_9_7,out_of_9_8,out_of_9_9,out_of_9_10,out_of_9_11,out_of_9_12,out_of_9_13,out_of_9_14,out_of_9_15,out_of_9_16,out_of_9_17,out_of_9_18,out_of_9_19,out_of_9_20,out_of_9_21,out_of_9_22,out_of_9_23,out_of_9_24,out_of_9_25,out_of_9_26,out_of_10_0,out_of_10_1,out_of_10_2,out_of_10_3,out_of_10_4,out_of_10_5,out_of_10_6,out_of_10_7,out_of_10_8,out_of_10_9,out_of_10_10,out_of_10_11,out_of_10_12,out_of_10_13,out_of_10_14,out_of_10_15,out_of_10_16,out_of_10_17,out_of_10_18,out_of_10_19,out_of_10_20,out_of_10_21,out_of_10_22,out_of_10_23,out_of_10_24,out_of_10_25,out_of_10_26,out_of_11_0,out_of_11_1,out_of_11_2,out_of_11_3,out_of_11_4,out_of_11_5,out_of_11_6,out_of_11_7,out_of_11_8,out_of_11_9,out_of_11_10,out_of_11_11,out_of_11_12,out_of_11_13,out_of_11_14,out_of_11_15,out_of_11_16,out_of_11_17,out_of_11_18,out_of_11_19,out_of_11_20,out_of_11_21,out_of_11_22,out_of_11_23,out_of_11_24,out_of_11_25,out_of_11_26,out_of_12_0,out_of_12_1,out_of_12_2,out_of_12_3,out_of_12_4,out_of_12_5,out_of_12_6,out_of_12_7,out_of_12_8,out_of_12_9,out_of_12_10,out_of_12_11,out_of_12_12,out_of_12_13,out_of_12_14,out_of_12_15,out_of_12_16,out_of_12_17,out_of_12_18,out_of_12_19,out_of_12_20,out_of_12_21,out_of_12_22,out_of_12_23,out_of_12_24,out_of_12_25,out_of_12_26,out_of_13_0,out_of_13_1,out_of_13_2,out_of_13_3,out_of_13_4,out_of_13_5,out_of_13_6,out_of_13_7,out_of_13_8,out_of_13_9,out_of_13_10,out_of_13_11,out_of_13_12,out_of_13_13,out_of_13_14,out_of_13_15,out_of_13_16,out_of_13_17,out_of_13_18,out_of_13_19,out_of_13_20,out_of_13_21,out_of_13_22,out_of_13_23,out_of_13_24,out_of_13_25,out_of_13_26,out_of_14_0,out_of_14_1,out_of_14_2,out_of_14_3,out_of_14_4,out_of_14_5,out_of_14_6,out_of_14_7,out_of_14_8,out_of_14_9,out_of_14_10,out_of_14_11,out_of_14_12,out_of_14_13,out_of_14_14,out_of_14_15,out_of_14_16,out_of_14_17,out_of_14_18,out_of_14_19,out_of_14_20,out_of_14_21,out_of_14_22,out_of_14_23,out_of_14_24,out_of_14_25,out_of_14_26,out_of_15_0,out_of_15_1,out_of_15_2,out_of_15_3,out_of_15_4,out_of_15_5,out_of_15_6,out_of_15_7,out_of_15_8,out_of_15_9,out_of_15_10,out_of_15_11,out_of_15_12,out_of_15_13,out_of_15_14,out_of_15_15,out_of_15_16,out_of_15_17,out_of_15_18,out_of_15_19,out_of_15_20,out_of_15_21,out_of_15_22,out_of_15_23,out_of_15_24,out_of_15_25,out_of_15_26;

reg [4:0] counter; // 27 cases, 27 differents sets of outputs all vertical.

//--------------------------------- Shift Register Horizontal -----------------------------//

register #(16) cell_0_0(clock, reset, enable, in_26, out_of_0_0);
register #(16) cell_0_1(clock, reset, enable, in_25, out_of_0_1);
register #(16) cell_0_2(clock, reset, enable, in_24, out_of_0_2);
register #(16) cell_0_3(clock, reset, enable, in_23, out_of_0_3);
register #(16) cell_0_4(clock, reset, enable, in_22, out_of_0_4);
register #(16) cell_0_5(clock, reset, enable, in_21, out_of_0_5);
register #(16) cell_0_6(clock, reset, enable, in_20, out_of_0_6);
register #(16) cell_0_7(clock, reset, enable, in_19, out_of_0_7);
register #(16) cell_0_8(clock, reset, enable, in_18, out_of_0_8);
register #(16) cell_0_9(clock, reset, enable, in_17, out_of_0_9);
register #(16) cell_0_10(clock, reset, enable, in_16, out_of_0_10);
register #(16) cell_0_11(clock, reset, enable, in_15, out_of_0_11);
register #(16) cell_0_12(clock, reset, enable, in_14, out_of_0_12);
register #(16) cell_0_13(clock, reset, enable, in_13, out_of_0_13);
register #(16) cell_0_14(clock, reset, enable, in_12, out_of_0_14);
register #(16) cell_0_15(clock, reset, enable, in_11, out_of_0_15);
register #(16) cell_0_16(clock, reset, enable, in_10, out_of_0_16);
register #(16) cell_0_17(clock, reset, enable, in_9, out_of_0_17);
register #(16) cell_0_18(clock, reset, enable, in_8, out_of_0_18);
register #(16) cell_0_19(clock, reset, enable, in_7, out_of_0_19);
register #(16) cell_0_20(clock, reset, enable, in_6, out_of_0_20);
register #(16) cell_0_21(clock, reset, enable, in_5, out_of_0_21);
register #(16) cell_0_22(clock, reset, enable, in_4, out_of_0_22);
register #(16) cell_0_23(clock, reset, enable, in_3, out_of_0_23);
register #(16) cell_0_24(clock, reset, enable, in_2, out_of_0_24);
register #(16) cell_0_25(clock, reset, enable, in_1, out_of_0_25);
register #(16) cell_0_26(clock, reset, enable, in_0, out_of_0_26);

register #(16) cell_1_0(clock, reset, enable, out_of_0_0, out_of_1_0);
register #(16) cell_1_1(clock, reset, enable, out_of_0_1, out_of_1_1);
register #(16) cell_1_2(clock, reset, enable, out_of_0_2, out_of_1_2);
register #(16) cell_1_3(clock, reset, enable, out_of_0_3, out_of_1_3);
register #(16) cell_1_4(clock, reset, enable, out_of_0_4, out_of_1_4);
register #(16) cell_1_5(clock, reset, enable, out_of_0_5, out_of_1_5);
register #(16) cell_1_6(clock, reset, enable, out_of_0_6, out_of_1_6);
register #(16) cell_1_7(clock, reset, enable, out_of_0_7, out_of_1_7);
register #(16) cell_1_8(clock, reset, enable, out_of_0_8, out_of_1_8);
register #(16) cell_1_9(clock, reset, enable, out_of_0_9, out_of_1_9);
register #(16) cell_1_10(clock, reset, enable, out_of_0_10, out_of_1_10);
register #(16) cell_1_11(clock, reset, enable,  out_of_0_11, out_of_1_11);
register #(16) cell_1_12(clock, reset, enable,  out_of_0_12, out_of_1_12);
register #(16) cell_1_13(clock, reset, enable,  out_of_0_13, out_of_1_13);
register #(16) cell_1_14(clock, reset, enable,  out_of_0_14, out_of_1_14);
register #(16) cell_1_15(clock, reset, enable,  out_of_0_15, out_of_1_15);
register #(16) cell_1_16(clock, reset, enable,  out_of_0_16, out_of_1_16);
register #(16) cell_1_17(clock, reset, enable,  out_of_0_17, out_of_1_17);
register #(16) cell_1_18(clock, reset, enable,  out_of_0_18, out_of_1_18);
register #(16) cell_1_19(clock, reset, enable,  out_of_0_19, out_of_1_19);
register #(16) cell_1_20(clock, reset, enable,  out_of_0_20, out_of_1_20);
register #(16) cell_1_21(clock, reset, enable,  out_of_0_21, out_of_1_21);
register #(16) cell_1_22(clock, reset, enable,  out_of_0_22, out_of_1_22);
register #(16) cell_1_23(clock, reset, enable,  out_of_0_23, out_of_1_23);
register #(16) cell_1_24(clock, reset, enable,  out_of_0_24, out_of_1_24);
register #(16) cell_1_25(clock, reset, enable,  out_of_0_25, out_of_1_25);
register #(16) cell_1_26(clock, reset, enable,  out_of_0_26, out_of_1_26);

register #(16) cell_2_0(clock, reset, enable,   out_of_1_0,  out_of_2_0);
register #(16) cell_2_1(clock, reset, enable,   out_of_1_1,  out_of_2_1);
register #(16) cell_2_2(clock, reset, enable,   out_of_1_2,  out_of_2_2);
register #(16) cell_2_3(clock, reset, enable,   out_of_1_3,  out_of_2_3);
register #(16) cell_2_4(clock, reset, enable,   out_of_1_4,  out_of_2_4);
register #(16) cell_2_5(clock, reset, enable,   out_of_1_5,  out_of_2_5);
register #(16) cell_2_6(clock, reset, enable,   out_of_1_6,  out_of_2_6);
register #(16) cell_2_7(clock, reset, enable,   out_of_1_7,  out_of_2_7);
register #(16) cell_2_8(clock, reset, enable,   out_of_1_8,  out_of_2_8);
register #(16) cell_2_9(clock, reset, enable,   out_of_1_9,  out_of_2_9);
register #(16) cell_2_10(clock, reset, enable,  out_of_1_10, out_of_2_10);
register #(16) cell_2_11(clock, reset, enable,  out_of_1_11, out_of_2_11);
register #(16) cell_2_12(clock, reset, enable,  out_of_1_12, out_of_2_12);
register #(16) cell_2_13(clock, reset, enable,  out_of_1_13, out_of_2_13);
register #(16) cell_2_14(clock, reset, enable,  out_of_1_14, out_of_2_14);
register #(16) cell_2_15(clock, reset, enable,  out_of_1_15, out_of_2_15);
register #(16) cell_2_16(clock, reset, enable,  out_of_1_16, out_of_2_16);
register #(16) cell_2_17(clock, reset, enable,  out_of_1_17, out_of_2_17);
register #(16) cell_2_18(clock, reset, enable,  out_of_1_18, out_of_2_18);
register #(16) cell_2_19(clock, reset, enable,  out_of_1_19, out_of_2_19);
register #(16) cell_2_20(clock, reset, enable,  out_of_1_20, out_of_2_20);
register #(16) cell_2_21(clock, reset, enable,  out_of_1_21, out_of_2_21);
register #(16) cell_2_22(clock, reset, enable,  out_of_1_22, out_of_2_22);
register #(16) cell_2_23(clock, reset, enable,  out_of_1_23, out_of_2_23);
register #(16) cell_2_24(clock, reset, enable,  out_of_1_24, out_of_2_24);
register #(16) cell_2_25(clock, reset, enable,  out_of_1_25, out_of_2_25);
register #(16) cell_2_26(clock, reset, enable,  out_of_1_26, out_of_2_26);

register #(16) cell_3_0(clock, reset, enable,   out_of_2_0,  out_of_3_0);
register #(16) cell_3_1(clock, reset, enable,   out_of_2_1,  out_of_3_1);
register #(16) cell_3_2(clock, reset, enable,   out_of_2_2,  out_of_3_2);
register #(16) cell_3_3(clock, reset, enable,   out_of_2_3,  out_of_3_3);
register #(16) cell_3_4(clock, reset, enable,   out_of_2_4,  out_of_3_4);
register #(16) cell_3_5(clock, reset, enable,   out_of_2_5,  out_of_3_5);
register #(16) cell_3_6(clock, reset, enable,   out_of_2_6,  out_of_3_6);
register #(16) cell_3_7(clock, reset, enable,   out_of_2_7,  out_of_3_7);
register #(16) cell_3_8(clock, reset, enable,   out_of_2_8,  out_of_3_8);
register #(16) cell_3_9(clock, reset, enable,   out_of_2_9,  out_of_3_9);
register #(16) cell_3_10(clock, reset, enable,  out_of_2_10, out_of_3_10);
register #(16) cell_3_11(clock, reset, enable,  out_of_2_11, out_of_3_11);
register #(16) cell_3_12(clock, reset, enable,  out_of_2_12, out_of_3_12);
register #(16) cell_3_13(clock, reset, enable,  out_of_2_13, out_of_3_13);
register #(16) cell_3_14(clock, reset, enable,  out_of_2_14, out_of_3_14);
register #(16) cell_3_15(clock, reset, enable,  out_of_2_15, out_of_3_15);
register #(16) cell_3_16(clock, reset, enable,  out_of_2_16, out_of_3_16);
register #(16) cell_3_17(clock, reset, enable,  out_of_2_17, out_of_3_17);
register #(16) cell_3_18(clock, reset, enable,  out_of_2_18, out_of_3_18);
register #(16) cell_3_19(clock, reset, enable,  out_of_2_19, out_of_3_19);
register #(16) cell_3_20(clock, reset, enable,  out_of_2_20, out_of_3_20);
register #(16) cell_3_21(clock, reset, enable,  out_of_2_21, out_of_3_21);
register #(16) cell_3_22(clock, reset, enable,  out_of_2_22, out_of_3_22);
register #(16) cell_3_23(clock, reset, enable,  out_of_2_23, out_of_3_23);
register #(16) cell_3_24(clock, reset, enable,  out_of_2_24, out_of_3_24);
register #(16) cell_3_25(clock, reset, enable,  out_of_2_25, out_of_3_25);
register #(16) cell_3_26(clock, reset, enable,  out_of_2_26, out_of_3_26);

register #(16) cell_4_0(clock, reset, enable,   out_of_3_0,  out_of_4_0);
register #(16) cell_4_1(clock, reset, enable,   out_of_3_1,  out_of_4_1);
register #(16) cell_4_2(clock, reset, enable,   out_of_3_2,  out_of_4_2);
register #(16) cell_4_3(clock, reset, enable,   out_of_3_3,  out_of_4_3);
register #(16) cell_4_4(clock, reset, enable,   out_of_3_4,  out_of_4_4);
register #(16) cell_4_5(clock, reset, enable,   out_of_3_5,  out_of_4_5);
register #(16) cell_4_6(clock, reset, enable,   out_of_3_6,  out_of_4_6);
register #(16) cell_4_7(clock, reset, enable,   out_of_3_7,  out_of_4_7);
register #(16) cell_4_8(clock, reset, enable,   out_of_3_8,  out_of_4_8);
register #(16) cell_4_9(clock, reset, enable,   out_of_3_9,  out_of_4_9);
register #(16) cell_4_10(clock, reset, enable,  out_of_3_10, out_of_4_10);
register #(16) cell_4_11(clock, reset, enable,  out_of_3_11, out_of_4_11);
register #(16) cell_4_12(clock, reset, enable,  out_of_3_12, out_of_4_12);
register #(16) cell_4_13(clock, reset, enable,  out_of_3_13, out_of_4_13);
register #(16) cell_4_14(clock, reset, enable,  out_of_3_14, out_of_4_14);
register #(16) cell_4_15(clock, reset, enable,  out_of_3_15, out_of_4_15);
register #(16) cell_4_16(clock, reset, enable,  out_of_3_16, out_of_4_16);
register #(16) cell_4_17(clock, reset, enable,  out_of_3_17, out_of_4_17);
register #(16) cell_4_18(clock, reset, enable,  out_of_3_18, out_of_4_18);
register #(16) cell_4_19(clock, reset, enable,  out_of_3_19, out_of_4_19);
register #(16) cell_4_20(clock, reset, enable,  out_of_3_20, out_of_4_20);
register #(16) cell_4_21(clock, reset, enable,  out_of_3_21, out_of_4_21);
register #(16) cell_4_22(clock, reset, enable,  out_of_3_22, out_of_4_22);
register #(16) cell_4_23(clock, reset, enable,  out_of_3_23, out_of_4_23);
register #(16) cell_4_24(clock, reset, enable,  out_of_3_24, out_of_4_24);
register #(16) cell_4_25(clock, reset, enable,  out_of_3_25, out_of_4_25);
register #(16) cell_4_26(clock, reset, enable,  out_of_3_26, out_of_4_26);

register #(16) cell_5_0(clock, reset, enable,   out_of_4_0,  out_of_5_0);
register #(16) cell_5_1(clock, reset, enable,   out_of_4_1,  out_of_5_1);
register #(16) cell_5_2(clock, reset, enable,   out_of_4_2,  out_of_5_2);
register #(16) cell_5_3(clock, reset, enable,   out_of_4_3,  out_of_5_3);
register #(16) cell_5_4(clock, reset, enable,   out_of_4_4,  out_of_5_4);
register #(16) cell_5_5(clock, reset, enable,   out_of_4_5,  out_of_5_5);
register #(16) cell_5_6(clock, reset, enable,   out_of_4_6,  out_of_5_6);
register #(16) cell_5_7(clock, reset, enable,   out_of_4_7,  out_of_5_7);
register #(16) cell_5_8(clock, reset, enable,   out_of_4_8,  out_of_5_8);
register #(16) cell_5_9(clock, reset, enable,   out_of_4_9,  out_of_5_9);
register #(16) cell_5_10(clock, reset, enable,  out_of_4_10, out_of_5_10);
register #(16) cell_5_11(clock, reset, enable,  out_of_4_11, out_of_5_11);
register #(16) cell_5_12(clock, reset, enable,  out_of_4_12, out_of_5_12);
register #(16) cell_5_13(clock, reset, enable,  out_of_4_13, out_of_5_13);
register #(16) cell_5_14(clock, reset, enable,  out_of_4_14, out_of_5_14);
register #(16) cell_5_15(clock, reset, enable,  out_of_4_15, out_of_5_15);
register #(16) cell_5_16(clock, reset, enable,  out_of_4_16, out_of_5_16);
register #(16) cell_5_17(clock, reset, enable,  out_of_4_17, out_of_5_17);
register #(16) cell_5_18(clock, reset, enable,  out_of_4_18, out_of_5_18);
register #(16) cell_5_19(clock, reset, enable,  out_of_4_19, out_of_5_19);
register #(16) cell_5_20(clock, reset, enable,  out_of_4_20, out_of_5_20);
register #(16) cell_5_21(clock, reset, enable,  out_of_4_21, out_of_5_21);
register #(16) cell_5_22(clock, reset, enable,  out_of_4_22, out_of_5_22);
register #(16) cell_5_23(clock, reset, enable,  out_of_4_23, out_of_5_23);
register #(16) cell_5_24(clock, reset, enable,  out_of_4_24, out_of_5_24);
register #(16) cell_5_25(clock, reset, enable,  out_of_4_25, out_of_5_25);
register #(16) cell_5_26(clock, reset, enable,  out_of_4_26, out_of_5_26);

register #(16) cell_6_0(clock, reset, enable,   out_of_5_0,  out_of_6_0);
register #(16) cell_6_1(clock, reset, enable,   out_of_5_1,  out_of_6_1);
register #(16) cell_6_2(clock, reset, enable,   out_of_5_2,  out_of_6_2);
register #(16) cell_6_3(clock, reset, enable,   out_of_5_3,  out_of_6_3);
register #(16) cell_6_4(clock, reset, enable,   out_of_5_4,  out_of_6_4);
register #(16) cell_6_5(clock, reset, enable,   out_of_5_5,  out_of_6_5);
register #(16) cell_6_6(clock, reset, enable,   out_of_5_6,  out_of_6_6);
register #(16) cell_6_7(clock, reset, enable,   out_of_5_7,  out_of_6_7);
register #(16) cell_6_8(clock, reset, enable,   out_of_5_8,  out_of_6_8);
register #(16) cell_6_9(clock, reset, enable,   out_of_5_9,  out_of_6_9);
register #(16) cell_6_10(clock, reset, enable,  out_of_5_10, out_of_6_10);
register #(16) cell_6_11(clock, reset, enable,  out_of_5_11, out_of_6_11);
register #(16) cell_6_12(clock, reset, enable,  out_of_5_12, out_of_6_12);
register #(16) cell_6_13(clock, reset, enable,  out_of_5_13, out_of_6_13);
register #(16) cell_6_14(clock, reset, enable,  out_of_5_14, out_of_6_14);
register #(16) cell_6_15(clock, reset, enable,  out_of_5_15, out_of_6_15);
register #(16) cell_6_16(clock, reset, enable,  out_of_5_16, out_of_6_16);
register #(16) cell_6_17(clock, reset, enable,  out_of_5_17, out_of_6_17);
register #(16) cell_6_18(clock, reset, enable,  out_of_5_18, out_of_6_18);
register #(16) cell_6_19(clock, reset, enable,  out_of_5_19, out_of_6_19);
register #(16) cell_6_20(clock, reset, enable,  out_of_5_20, out_of_6_20);
register #(16) cell_6_21(clock, reset, enable,  out_of_5_21, out_of_6_21);
register #(16) cell_6_22(clock, reset, enable,  out_of_5_22, out_of_6_22);
register #(16) cell_6_23(clock, reset, enable,  out_of_5_23, out_of_6_23);
register #(16) cell_6_24(clock, reset, enable,  out_of_5_24, out_of_6_24);
register #(16) cell_6_25(clock, reset, enable,  out_of_5_25, out_of_6_25);
register #(16) cell_6_26(clock, reset, enable,  out_of_5_26, out_of_6_26);

register #(16) cell_7_0(clock, reset, enable,   out_of_6_0,  out_of_7_0);
register #(16) cell_7_1(clock, reset, enable,   out_of_6_1,  out_of_7_1);
register #(16) cell_7_2(clock, reset, enable,   out_of_6_2,  out_of_7_2);
register #(16) cell_7_3(clock, reset, enable,   out_of_6_3,  out_of_7_3);
register #(16) cell_7_4(clock, reset, enable,   out_of_6_4,  out_of_7_4);
register #(16) cell_7_5(clock, reset, enable,   out_of_6_5,  out_of_7_5);
register #(16) cell_7_6(clock, reset, enable,   out_of_6_6,  out_of_7_6);
register #(16) cell_7_7(clock, reset, enable,   out_of_6_7,  out_of_7_7);
register #(16) cell_7_8(clock, reset, enable,   out_of_6_8,  out_of_7_8);
register #(16) cell_7_9(clock, reset, enable,   out_of_6_9,  out_of_7_9);
register #(16) cell_7_10(clock, reset, enable,  out_of_6_10, out_of_7_10);
register #(16) cell_7_11(clock, reset, enable,  out_of_6_11, out_of_7_11);
register #(16) cell_7_12(clock, reset, enable,  out_of_6_12, out_of_7_12);
register #(16) cell_7_13(clock, reset, enable,  out_of_6_13, out_of_7_13);
register #(16) cell_7_14(clock, reset, enable,  out_of_6_14, out_of_7_14);
register #(16) cell_7_15(clock, reset, enable,  out_of_6_15, out_of_7_15);
register #(16) cell_7_16(clock, reset, enable,  out_of_6_16, out_of_7_16);
register #(16) cell_7_17(clock, reset, enable,  out_of_6_17, out_of_7_17);
register #(16) cell_7_18(clock, reset, enable,  out_of_6_18, out_of_7_18);
register #(16) cell_7_19(clock, reset, enable,  out_of_6_19, out_of_7_19);
register #(16) cell_7_20(clock, reset, enable,  out_of_6_20, out_of_7_20);
register #(16) cell_7_21(clock, reset, enable,  out_of_6_21, out_of_7_21);
register #(16) cell_7_22(clock, reset, enable,  out_of_6_22, out_of_7_22);
register #(16) cell_7_23(clock, reset, enable,  out_of_6_23, out_of_7_23);
register #(16) cell_7_24(clock, reset, enable,  out_of_6_24, out_of_7_24);
register #(16) cell_7_25(clock, reset, enable,  out_of_6_25, out_of_7_25);
register #(16) cell_7_26(clock, reset, enable,  out_of_6_26, out_of_7_26);

register #(16) cell_8_0(clock, reset, enable,   out_of_7_0,  out_of_8_0);
register #(16) cell_8_1(clock, reset, enable,   out_of_7_1,  out_of_8_1);
register #(16) cell_8_2(clock, reset, enable,   out_of_7_2,  out_of_8_2);
register #(16) cell_8_3(clock, reset, enable,   out_of_7_3,  out_of_8_3);
register #(16) cell_8_4(clock, reset, enable,   out_of_7_4,  out_of_8_4);
register #(16) cell_8_5(clock, reset, enable,   out_of_7_5,  out_of_8_5);
register #(16) cell_8_6(clock, reset, enable,   out_of_7_6,  out_of_8_6);
register #(16) cell_8_7(clock, reset, enable,   out_of_7_7,  out_of_8_7);
register #(16) cell_8_8(clock, reset, enable,   out_of_7_8,  out_of_8_8);
register #(16) cell_8_9(clock, reset, enable,   out_of_7_9,  out_of_8_9);
register #(16) cell_8_10(clock, reset, enable,  out_of_7_10, out_of_8_10);
register #(16) cell_8_11(clock, reset, enable,  out_of_7_11, out_of_8_11);
register #(16) cell_8_12(clock, reset, enable,  out_of_7_12, out_of_8_12);
register #(16) cell_8_13(clock, reset, enable,  out_of_7_13, out_of_8_13);
register #(16) cell_8_14(clock, reset, enable,  out_of_7_14, out_of_8_14);
register #(16) cell_8_15(clock, reset, enable,  out_of_7_15, out_of_8_15);
register #(16) cell_8_16(clock, reset, enable,  out_of_7_16, out_of_8_16);
register #(16) cell_8_17(clock, reset, enable,  out_of_7_17, out_of_8_17);
register #(16) cell_8_18(clock, reset, enable,  out_of_7_18, out_of_8_18);
register #(16) cell_8_19(clock, reset, enable,  out_of_7_19, out_of_8_19);
register #(16) cell_8_20(clock, reset, enable,  out_of_7_20, out_of_8_20);
register #(16) cell_8_21(clock, reset, enable,  out_of_7_21, out_of_8_21);
register #(16) cell_8_22(clock, reset, enable,  out_of_7_22, out_of_8_22);
register #(16) cell_8_23(clock, reset, enable,  out_of_7_23, out_of_8_23);
register #(16) cell_8_24(clock, reset, enable,  out_of_7_24, out_of_8_24);
register #(16) cell_8_25(clock, reset, enable,  out_of_7_25, out_of_8_25);
register #(16) cell_8_26(clock, reset, enable,  out_of_7_26, out_of_8_26);

register #(16) cell_9_0(clock, reset, enable,   out_of_8_0,  out_of_9_0);
register #(16) cell_9_1(clock, reset, enable,   out_of_8_1,  out_of_9_1);
register #(16) cell_9_2(clock, reset, enable,   out_of_8_2,  out_of_9_2);
register #(16) cell_9_3(clock, reset, enable,   out_of_8_3,  out_of_9_3);
register #(16) cell_9_4(clock, reset, enable,   out_of_8_4,  out_of_9_4);
register #(16) cell_9_5(clock, reset, enable,   out_of_8_5,  out_of_9_5);
register #(16) cell_9_6(clock, reset, enable,   out_of_8_6,  out_of_9_6);
register #(16) cell_9_7(clock, reset, enable,   out_of_8_7,  out_of_9_7);
register #(16) cell_9_8(clock, reset, enable,   out_of_8_8,  out_of_9_8);
register #(16) cell_9_9(clock, reset, enable,   out_of_8_9,  out_of_9_9);
register #(16) cell_9_10(clock, reset, enable,  out_of_8_10, out_of_9_10);
register #(16) cell_9_11(clock, reset, enable,  out_of_8_11, out_of_9_11);
register #(16) cell_9_12(clock, reset, enable,  out_of_8_12, out_of_9_12);
register #(16) cell_9_13(clock, reset, enable,  out_of_8_13, out_of_9_13);
register #(16) cell_9_14(clock, reset, enable,  out_of_8_14, out_of_9_14);
register #(16) cell_9_15(clock, reset, enable,  out_of_8_15, out_of_9_15);
register #(16) cell_9_16(clock, reset, enable,  out_of_8_16, out_of_9_16);
register #(16) cell_9_17(clock, reset, enable,  out_of_8_17, out_of_9_17);
register #(16) cell_9_18(clock, reset, enable,  out_of_8_18, out_of_9_18);
register #(16) cell_9_19(clock, reset, enable,  out_of_8_19, out_of_9_19);
register #(16) cell_9_20(clock, reset, enable,  out_of_8_20, out_of_9_20);
register #(16) cell_9_21(clock, reset, enable,  out_of_8_21, out_of_9_21);
register #(16) cell_9_22(clock, reset, enable,  out_of_8_22, out_of_9_22);
register #(16) cell_9_23(clock, reset, enable,  out_of_8_23, out_of_9_23);
register #(16) cell_9_24(clock, reset, enable,  out_of_8_24, out_of_9_24);
register #(16) cell_9_25(clock, reset, enable,  out_of_8_25, out_of_9_25);
register #(16) cell_9_26(clock, reset, enable,  out_of_8_26, out_of_9_26);

register #(16) cell_10_0(clock, reset, enable,   out_of_9_0,  out_of_10_0);
register #(16) cell_10_1(clock, reset, enable,   out_of_9_1,  out_of_10_1);
register #(16) cell_10_2(clock, reset, enable,   out_of_9_2,  out_of_10_2);
register #(16) cell_10_3(clock, reset, enable,   out_of_9_3,  out_of_10_3);
register #(16) cell_10_4(clock, reset, enable,   out_of_9_4,  out_of_10_4);
register #(16) cell_10_5(clock, reset, enable,   out_of_9_5,  out_of_10_5);
register #(16) cell_10_6(clock, reset, enable,   out_of_9_6,  out_of_10_6);
register #(16) cell_10_7(clock, reset, enable,   out_of_9_7,  out_of_10_7);
register #(16) cell_10_8(clock, reset, enable,   out_of_9_8,  out_of_10_8);
register #(16) cell_10_9(clock, reset, enable,   out_of_9_9,  out_of_10_9);
register #(16) cell_10_10(clock, reset, enable,  out_of_9_10, out_of_10_10);
register #(16) cell_10_11(clock, reset, enable,  out_of_9_11, out_of_10_11);
register #(16) cell_10_12(clock, reset, enable,  out_of_9_12, out_of_10_12);
register #(16) cell_10_13(clock, reset, enable,  out_of_9_13, out_of_10_13);
register #(16) cell_10_14(clock, reset, enable,  out_of_9_14, out_of_10_14);
register #(16) cell_10_15(clock, reset, enable,  out_of_9_15, out_of_10_15);
register #(16) cell_10_16(clock, reset, enable,  out_of_9_16, out_of_10_16);
register #(16) cell_10_17(clock, reset, enable,  out_of_9_17, out_of_10_17);
register #(16) cell_10_18(clock, reset, enable,  out_of_9_18, out_of_10_18);
register #(16) cell_10_19(clock, reset, enable,  out_of_9_19, out_of_10_19);
register #(16) cell_10_20(clock, reset, enable,  out_of_9_20, out_of_10_20);
register #(16) cell_10_21(clock, reset, enable,  out_of_9_21, out_of_10_21);
register #(16) cell_10_22(clock, reset, enable,  out_of_9_22, out_of_10_22);
register #(16) cell_10_23(clock, reset, enable,  out_of_9_23, out_of_10_23);
register #(16) cell_10_24(clock, reset, enable,  out_of_9_24, out_of_10_24);
register #(16) cell_10_25(clock, reset, enable,  out_of_9_25, out_of_10_25);
register #(16) cell_10_26(clock, reset, enable,  out_of_9_26, out_of_10_26);

register #(16) cell_11_0(clock, reset, enable,   out_of_10_0,  out_of_11_0);
register #(16) cell_11_1(clock, reset, enable,   out_of_10_1,  out_of_11_1);
register #(16) cell_11_2(clock, reset, enable,   out_of_10_2,  out_of_11_2);
register #(16) cell_11_3(clock, reset, enable,   out_of_10_3,  out_of_11_3);
register #(16) cell_11_4(clock, reset, enable,   out_of_10_4,  out_of_11_4);
register #(16) cell_11_5(clock, reset, enable,   out_of_10_5,  out_of_11_5);
register #(16) cell_11_6(clock, reset, enable,   out_of_10_6,  out_of_11_6);
register #(16) cell_11_7(clock, reset, enable,   out_of_10_7,  out_of_11_7);
register #(16) cell_11_8(clock, reset, enable,   out_of_10_8,  out_of_11_8);
register #(16) cell_11_9(clock, reset, enable,   out_of_10_9,  out_of_11_9);
register #(16) cell_11_10(clock, reset, enable,  out_of_10_10, out_of_11_10);
register #(16) cell_11_11(clock, reset, enable,  out_of_10_11, out_of_11_11);
register #(16) cell_11_12(clock, reset, enable,  out_of_10_12, out_of_11_12);
register #(16) cell_11_13(clock, reset, enable,  out_of_10_13, out_of_11_13);
register #(16) cell_11_14(clock, reset, enable,  out_of_10_14, out_of_11_14);
register #(16) cell_11_15(clock, reset, enable,  out_of_10_15, out_of_11_15);
register #(16) cell_11_16(clock, reset, enable,  out_of_10_16, out_of_11_16);
register #(16) cell_11_17(clock, reset, enable,  out_of_10_17, out_of_11_17);
register #(16) cell_11_18(clock, reset, enable,  out_of_10_18, out_of_11_18);
register #(16) cell_11_19(clock, reset, enable,  out_of_10_19, out_of_11_19);
register #(16) cell_11_20(clock, reset, enable,  out_of_10_20, out_of_11_20);
register #(16) cell_11_21(clock, reset, enable,  out_of_10_21, out_of_11_21);
register #(16) cell_11_22(clock, reset, enable,  out_of_10_22, out_of_11_22);
register #(16) cell_11_23(clock, reset, enable,  out_of_10_23, out_of_11_23);
register #(16) cell_11_24(clock, reset, enable,  out_of_10_24, out_of_11_24);
register #(16) cell_11_25(clock, reset, enable,  out_of_10_25, out_of_11_25);
register #(16) cell_11_26(clock, reset, enable,  out_of_10_26, out_of_11_26);
register #(16) cell_12_0(clock, reset, enable,   out_of_11_0,  out_of_12_0);
register #(16) cell_12_1(clock, reset, enable,   out_of_11_1,  out_of_12_1);
register #(16) cell_12_2(clock, reset, enable,   out_of_11_2,  out_of_12_2);
register #(16) cell_12_3(clock, reset, enable,   out_of_11_3,  out_of_12_3);
register #(16) cell_12_4(clock, reset, enable,   out_of_11_4,  out_of_12_4);
register #(16) cell_12_5(clock, reset, enable,   out_of_11_5,  out_of_12_5);
register #(16) cell_12_6(clock, reset, enable,   out_of_11_6,  out_of_12_6);
register #(16) cell_12_7(clock, reset, enable,   out_of_11_7,  out_of_12_7);
register #(16) cell_12_8(clock, reset, enable,   out_of_11_8,  out_of_12_8);
register #(16) cell_12_9(clock, reset, enable,   out_of_11_9,  out_of_12_9);
register #(16) cell_12_10(clock, reset, enable,  out_of_11_10, out_of_12_10);
register #(16) cell_12_11(clock, reset, enable,  out_of_11_11, out_of_12_11);
register #(16) cell_12_12(clock, reset, enable,  out_of_11_12, out_of_12_12);
register #(16) cell_12_13(clock, reset, enable,  out_of_11_13, out_of_12_13);
register #(16) cell_12_14(clock, reset, enable,  out_of_11_14, out_of_12_14);
register #(16) cell_12_15(clock, reset, enable,  out_of_11_15, out_of_12_15);
register #(16) cell_12_16(clock, reset, enable,  out_of_11_16, out_of_12_16);
register #(16) cell_12_17(clock, reset, enable,  out_of_11_17, out_of_12_17);
register #(16) cell_12_18(clock, reset, enable,  out_of_11_18, out_of_12_18);
register #(16) cell_12_19(clock, reset, enable,  out_of_11_19, out_of_12_19);
register #(16) cell_12_20(clock, reset, enable,  out_of_11_20, out_of_12_20);
register #(16) cell_12_21(clock, reset, enable,  out_of_11_21, out_of_12_21);
register #(16) cell_12_22(clock, reset, enable,  out_of_11_22, out_of_12_22);
register #(16) cell_12_23(clock, reset, enable,  out_of_11_23, out_of_12_23);
register #(16) cell_12_24(clock, reset, enable,  out_of_11_24, out_of_12_24);
register #(16) cell_12_25(clock, reset, enable,  out_of_11_25, out_of_12_25);
register #(16) cell_12_26(clock, reset, enable,  out_of_11_26, out_of_12_26);
register #(16) cell_13_0(clock, reset, enable,   out_of_12_0,  out_of_13_0);
register #(16) cell_13_1(clock, reset, enable,   out_of_12_1,  out_of_13_1);
register #(16) cell_13_2(clock, reset, enable,   out_of_12_2,  out_of_13_2);
register #(16) cell_13_3(clock, reset, enable,   out_of_12_3,  out_of_13_3);
register #(16) cell_13_4(clock, reset, enable,   out_of_12_4,  out_of_13_4);
register #(16) cell_13_5(clock, reset, enable,   out_of_12_5,  out_of_13_5);
register #(16) cell_13_6(clock, reset, enable,   out_of_12_6,  out_of_13_6);
register #(16) cell_13_7(clock, reset, enable,   out_of_12_7,  out_of_13_7);
register #(16) cell_13_8(clock, reset, enable,   out_of_12_8,  out_of_13_8);
register #(16) cell_13_9(clock, reset, enable,   out_of_12_9,  out_of_13_9);
register #(16) cell_13_10(clock, reset, enable,  out_of_12_10, out_of_13_10);
register #(16) cell_13_11(clock, reset, enable,  out_of_12_11, out_of_13_11);
register #(16) cell_13_12(clock, reset, enable,  out_of_12_12, out_of_13_12);
register #(16) cell_13_13(clock, reset, enable,  out_of_12_13, out_of_13_13);
register #(16) cell_13_14(clock, reset, enable,  out_of_12_14, out_of_13_14);
register #(16) cell_13_15(clock, reset, enable,  out_of_12_15, out_of_13_15);
register #(16) cell_13_16(clock, reset, enable,  out_of_12_16, out_of_13_16);
register #(16) cell_13_17(clock, reset, enable,  out_of_12_17, out_of_13_17);
register #(16) cell_13_18(clock, reset, enable,  out_of_12_18, out_of_13_18);
register #(16) cell_13_19(clock, reset, enable,  out_of_12_19, out_of_13_19);
register #(16) cell_13_20(clock, reset, enable,  out_of_12_20, out_of_13_20);
register #(16) cell_13_21(clock, reset, enable,  out_of_12_21, out_of_13_21);
register #(16) cell_13_22(clock, reset, enable,  out_of_12_22, out_of_13_22);
register #(16) cell_13_23(clock, reset, enable,  out_of_12_23, out_of_13_23);
register #(16) cell_13_24(clock, reset, enable,  out_of_12_24, out_of_13_24);
register #(16) cell_13_25(clock, reset, enable,  out_of_12_25, out_of_13_25);
register #(16) cell_13_26(clock, reset, enable,  out_of_12_26, out_of_13_26);
register #(16) cell_14_0(clock, reset, enable,   out_of_13_0,   out_of_14_0);
register #(16) cell_14_1(clock, reset, enable,   out_of_13_1,   out_of_14_1);
register #(16) cell_14_2(clock, reset, enable,   out_of_13_2,   out_of_14_2);
register #(16) cell_14_3(clock, reset, enable,   out_of_13_3,   out_of_14_3);
register #(16) cell_14_4(clock, reset, enable,   out_of_13_4,   out_of_14_4);
register #(16) cell_14_5(clock, reset, enable,   out_of_13_5,   out_of_14_5);
register #(16) cell_14_6(clock, reset, enable,   out_of_13_6,   out_of_14_6);
register #(16) cell_14_7(clock, reset, enable,   out_of_13_7,   out_of_14_7);
register #(16) cell_14_8(clock, reset, enable,   out_of_13_8,   out_of_14_8);
register #(16) cell_14_9(clock, reset, enable,   out_of_13_9,   out_of_14_9);
register #(16) cell_14_10(clock, reset, enable,  out_of_13_10,  out_of_14_10);
register #(16) cell_14_11(clock, reset, enable,  out_of_13_11,  out_of_14_11);
register #(16) cell_14_12(clock, reset, enable,  out_of_13_12,  out_of_14_12);
register #(16) cell_14_13(clock, reset, enable,  out_of_13_13,  out_of_14_13);
register #(16) cell_14_14(clock, reset, enable,  out_of_13_14,  out_of_14_14);
register #(16) cell_14_15(clock, reset, enable,  out_of_13_15,  out_of_14_15);
register #(16) cell_14_16(clock, reset, enable,  out_of_13_16,  out_of_14_16);
register #(16) cell_14_17(clock, reset, enable,  out_of_13_17,  out_of_14_17);
register #(16) cell_14_18(clock, reset, enable,  out_of_13_18,  out_of_14_18);
register #(16) cell_14_19(clock, reset, enable,  out_of_13_19,  out_of_14_19);
register #(16) cell_14_20(clock, reset, enable,  out_of_13_20,  out_of_14_20);
register #(16) cell_14_21(clock, reset, enable,  out_of_13_21,  out_of_14_21);
register #(16) cell_14_22(clock, reset, enable,  out_of_13_22,  out_of_14_22);
register #(16) cell_14_23(clock, reset, enable,  out_of_13_23,  out_of_14_23);
register #(16) cell_14_24(clock, reset, enable,  out_of_13_24,  out_of_14_24);
register #(16) cell_14_25(clock, reset, enable,  out_of_13_25,  out_of_14_25);
register #(16) cell_14_26(clock, reset, enable,  out_of_13_26,  out_of_14_26);
register #(16) cell_15_0(clock, reset, enable,   out_of_14_0,   out_of_15_0);
register #(16) cell_15_1(clock, reset, enable,   out_of_14_1,   out_of_15_1);
register #(16) cell_15_2(clock, reset, enable,   out_of_14_2,   out_of_15_2);
register #(16) cell_15_3(clock, reset, enable,   out_of_14_3,   out_of_15_3);
register #(16) cell_15_4(clock, reset, enable,   out_of_14_4,   out_of_15_4);
register #(16) cell_15_5(clock, reset, enable,   out_of_14_5,   out_of_15_5);
register #(16) cell_15_6(clock, reset, enable,   out_of_14_6,   out_of_15_6);
register #(16) cell_15_7(clock, reset, enable,   out_of_14_7,   out_of_15_7);
register #(16) cell_15_8(clock, reset, enable,   out_of_14_8,   out_of_15_8);
register #(16) cell_15_9(clock, reset, enable,   out_of_14_9,   out_of_15_9);
register #(16) cell_15_10(clock, reset, enable,  out_of_14_10,  out_of_15_10);
register #(16) cell_15_11(clock, reset, enable,  out_of_14_11,  out_of_15_11);
register #(16) cell_15_12(clock, reset, enable,  out_of_14_12,  out_of_15_12);
register #(16) cell_15_13(clock, reset, enable,  out_of_14_13,  out_of_15_13);
register #(16) cell_15_14(clock, reset, enable,  out_of_14_14,  out_of_15_14);
register #(16) cell_15_15(clock, reset, enable,  out_of_14_15,  out_of_15_15);
register #(16) cell_15_16(clock, reset, enable,  out_of_14_16,  out_of_15_16);
register #(16) cell_15_17(clock, reset, enable,  out_of_14_17,  out_of_15_17);
register #(16) cell_15_18(clock, reset, enable,  out_of_14_18,  out_of_15_18);
register #(16) cell_15_19(clock, reset, enable,  out_of_14_19,  out_of_15_19);
register #(16) cell_15_20(clock, reset, enable,  out_of_14_20,  out_of_15_20);
register #(16) cell_15_21(clock, reset, enable,  out_of_14_21,  out_of_15_21);
register #(16) cell_15_22(clock, reset, enable,  out_of_14_22,  out_of_15_22);
register #(16) cell_15_23(clock, reset, enable,  out_of_14_23,  out_of_15_23);
register #(16) cell_15_24(clock, reset, enable,  out_of_14_24,  out_of_15_24);
register #(16) cell_15_25(clock, reset, enable,  out_of_14_25,  out_of_15_25);
register #(16) cell_15_26(clock, reset, enable,  out_of_14_26,  out_of_15_26);

always @(posedge clock or posedge reset) begin 
 	if (reset) begin
 		counter <= 0;
 	end
 	else if (enable) begin
 		counter <= 0;
 	end
 	else if (enable_read) begin
 		counter <= counter +1;
 	end
 	else begin
 		counter <= 1;
 	end
 end

always @ (posedge clock )
case (counter)
  5'b00000 : 
	begin
	out_0 <=  0; 
	out_1 <=  0; 
	out_2 <=  0; 
	out_3 <=  0; 
	out_4 <=  0; 
	out_5 <=  0; 
	out_6 <=  0; 
	out_7 <=  0; 
	out_8 <=  0; 
	out_9 <=  0; 
	out_10 <= 0;
	out_11 <= 0;
	out_12 <= 0;
	out_13 <= 0;
	out_14 <= 0;
	out_15 <= 0;
	end

  5'b00001 : 	
	begin
	out_0 <=   out_of_0_26; 
	out_1 <=   out_of_1_26; 
	out_2 <=   out_of_2_26; 
	out_3 <=   out_of_3_26; 
	out_4 <=   out_of_4_26; 
	out_5 <=   out_of_5_26; 
	out_6 <=   out_of_6_26; 
	out_7 <=   out_of_7_26; 
	out_8 <=   out_of_8_26; 
	out_9 <=   out_of_9_26; 
	out_10 <= out_of_10_26;
	out_11 <= out_of_11_26;
	out_12 <= out_of_12_26;
	out_13 <= out_of_13_26;
	out_14 <= out_of_14_26;
	out_15 <= out_of_15_26;
	end

  5'b00010 : 	
	begin
	out_0 <=   out_of_0_25; 
	out_1 <=   out_of_1_25; 
	out_2 <=   out_of_2_25; 
	out_3 <=   out_of_3_25; 
	out_4 <=   out_of_4_25; 
	out_5 <=   out_of_5_25; 
	out_6 <=   out_of_6_25; 
	out_7 <=   out_of_7_25; 
	out_8 <=   out_of_8_25; 
	out_9 <=   out_of_9_25; 
	out_10 <= out_of_10_25;
	out_11 <= out_of_11_25;
	out_12 <= out_of_12_25;
	out_13 <= out_of_13_25;
	out_14 <= out_of_14_25;
	out_15 <= out_of_15_25;
	end
  5'b00011 : 	
	begin
	out_0 <=   out_of_0_24; 
	out_1 <=   out_of_1_24; 
	out_2 <=   out_of_2_24; 
	out_3 <=   out_of_3_24; 
	out_4 <=   out_of_4_24; 
	out_5 <=   out_of_5_24; 
	out_6 <=   out_of_6_24; 
	out_7 <=   out_of_7_24; 
	out_8 <=   out_of_8_24; 
	out_9 <=   out_of_9_24; 
	out_10 <= out_of_10_24;
	out_11 <= out_of_11_24;
	out_12 <= out_of_12_24;
	out_13 <= out_of_13_24;
	out_14 <= out_of_14_24;
	out_15 <= out_of_15_24;
	end
  5'b00100 : 	
	begin
	out_0 <=   out_of_0_23; 
	out_1 <=   out_of_1_23; 
	out_2 <=   out_of_2_23; 
	out_3 <=   out_of_3_23; 
	out_4 <=   out_of_4_23; 
	out_5 <=   out_of_5_23; 
	out_6 <=   out_of_6_23; 
	out_7 <=   out_of_7_23; 
	out_8 <=   out_of_8_23; 
	out_9 <=   out_of_9_23; 
	out_10 <= out_of_10_23;
	out_11 <= out_of_11_23;
	out_12 <= out_of_12_23;
	out_13 <= out_of_13_23;
	out_14 <= out_of_14_23;
	out_15 <= out_of_15_23;
	end
  5'b00101 : 	
	begin
	out_0 <=   out_of_0_22; 
	out_1 <=   out_of_1_22; 
	out_2 <=   out_of_2_22; 
	out_3 <=   out_of_3_22; 
	out_4 <=   out_of_4_22; 
	out_5 <=   out_of_5_22; 
	out_6 <=   out_of_6_22; 
	out_7 <=   out_of_7_22; 
	out_8 <=   out_of_8_22; 
	out_9 <=   out_of_9_22; 
	out_10 <= out_of_10_22;
	out_11 <= out_of_11_22;
	out_12 <= out_of_12_22;
	out_13 <= out_of_13_22;
	out_14 <= out_of_14_22;
	out_15 <= out_of_15_22;
	end
  5'b00110 : 	
	begin
	out_0 <=   out_of_0_21; 
	out_1 <=   out_of_1_21; 
	out_2 <=   out_of_2_21; 
	out_3 <=   out_of_3_21; 
	out_4 <=   out_of_4_21; 
	out_5 <=   out_of_5_21; 
	out_6 <=   out_of_6_21; 
	out_7 <=   out_of_7_21; 
	out_8 <=   out_of_8_21; 
	out_9 <=   out_of_9_21; 
	out_10 <= out_of_10_21;
	out_11 <= out_of_11_21;
	out_12 <= out_of_12_21;
	out_13 <= out_of_13_21;
	out_14 <= out_of_14_21;
	out_15 <= out_of_15_21;
	end
  5'b00111 : 	
	begin
	out_0 <=   out_of_0_20; 
	out_1 <=   out_of_1_20; 
	out_2 <=   out_of_2_20; 
	out_3 <=   out_of_3_20; 
	out_4 <=   out_of_4_20; 
	out_5 <=   out_of_5_20; 
	out_6 <=   out_of_6_20; 
	out_7 <=   out_of_7_20; 
	out_8 <=   out_of_8_20; 
	out_9 <=   out_of_9_20; 
	out_10 <= out_of_10_20;
	out_11 <= out_of_11_20;
	out_12 <= out_of_12_20;
	out_13 <= out_of_13_20;
	out_14 <= out_of_14_20;
	out_15 <= out_of_15_20;
	end



  5'b01000 : 
	begin
	out_0 <=   out_of_0_19; 
	out_1 <=   out_of_1_19; 
	out_2 <=   out_of_2_19; 
	out_3 <=   out_of_3_19; 
	out_4 <=   out_of_4_19; 
	out_5 <=   out_of_5_19; 
	out_6 <=   out_of_6_19; 
	out_7 <=   out_of_7_19; 
	out_8 <=   out_of_8_19; 
	out_9 <=   out_of_9_19; 
	out_10 <= out_of_10_19;
	out_11 <= out_of_11_19;
	out_12 <= out_of_12_19;
	out_13 <= out_of_13_19;
	out_14 <= out_of_14_19;
	out_15 <= out_of_15_19;
	end

  5'b01001 : 	
	begin
	out_0 <=   out_of_0_18; 
	out_1 <=   out_of_1_18; 
	out_2 <=   out_of_2_18; 
	out_3 <=   out_of_3_18; 
	out_4 <=   out_of_4_18; 
	out_5 <=   out_of_5_18; 
	out_6 <=   out_of_6_18; 
	out_7 <=   out_of_7_18; 
	out_8 <=   out_of_8_18; 
	out_9 <=   out_of_9_18; 
	out_10 <= out_of_10_18;
	out_11 <= out_of_11_18;
	out_12 <= out_of_12_18;
	out_13 <= out_of_13_18;
	out_14 <= out_of_14_18;
	out_15 <= out_of_15_18;
	end

  5'b01010 : 	
	begin
	out_0 <=   out_of_0_17; 
	out_1 <=   out_of_1_17; 
	out_2 <=   out_of_2_17; 
	out_3 <=   out_of_3_17; 
	out_4 <=   out_of_4_17; 
	out_5 <=   out_of_5_17; 
	out_6 <=   out_of_6_17; 
	out_7 <=   out_of_7_17; 
	out_8 <=   out_of_8_17; 
	out_9 <=   out_of_9_17; 
	out_10 <= out_of_10_17;
	out_11 <= out_of_11_17;
	out_12 <= out_of_12_17;
	out_13 <= out_of_13_17;
	out_14 <= out_of_14_17;
	out_15 <= out_of_15_17;
	end
  5'b01011 : 	
	begin
	out_0 <=   out_of_0_16; 
	out_1 <=   out_of_1_16; 
	out_2 <=   out_of_2_16; 
	out_3 <=   out_of_3_16; 
	out_4 <=   out_of_4_16; 
	out_5 <=   out_of_5_16; 
	out_6 <=   out_of_6_16; 
	out_7 <=   out_of_7_16; 
	out_8 <=   out_of_8_16; 
	out_9 <=   out_of_9_16; 
	out_10 <= out_of_10_16;
	out_11 <= out_of_11_16;
	out_12 <= out_of_12_16;
	out_13 <= out_of_13_16;
	out_14 <= out_of_14_16;
	out_15 <= out_of_15_16;
	end
  5'b01100 : 	
	begin
	out_0 <=   out_of_0_15; 
	out_1 <=   out_of_1_15; 
	out_2 <=   out_of_2_15; 
	out_3 <=   out_of_3_15; 
	out_4 <=   out_of_4_15; 
	out_5 <=   out_of_5_15; 
	out_6 <=   out_of_6_15; 
	out_7 <=   out_of_7_15; 
	out_8 <=   out_of_8_15; 
	out_9 <=   out_of_9_15; 
	out_10 <= out_of_10_15;
	out_11 <= out_of_11_15;
	out_12 <= out_of_12_15;
	out_13 <= out_of_13_15;
	out_14 <= out_of_14_15;
	out_15 <= out_of_15_15;
	end
  5'b01101 : 	
	begin
	out_0 <=   out_of_0_14; 
	out_1 <=   out_of_1_14; 
	out_2 <=   out_of_2_14; 
	out_3 <=   out_of_3_14; 
	out_4 <=   out_of_4_14; 
	out_5 <=   out_of_5_14; 
	out_6 <=   out_of_6_14; 
	out_7 <=   out_of_7_14; 
	out_8 <=   out_of_8_14; 
	out_9 <=   out_of_9_14; 
	out_10 <= out_of_10_14;
	out_11 <= out_of_11_14;
	out_12 <= out_of_12_14;
	out_13 <= out_of_13_14;
	out_14 <= out_of_14_14;
	out_15 <= out_of_15_14;
	end
  5'b01110 : 	
	begin
	out_0 <=   out_of_0_13; 
	out_1 <=   out_of_1_13; 
	out_2 <=   out_of_2_13; 
	out_3 <=   out_of_3_13; 
	out_4 <=   out_of_4_13; 
	out_5 <=   out_of_5_13; 
	out_6 <=   out_of_6_13; 
	out_7 <=   out_of_7_13; 
	out_8 <=   out_of_8_13; 
	out_9 <=   out_of_9_13; 
	out_10 <= out_of_10_13;
	out_11 <= out_of_11_13;
	out_12 <= out_of_12_13;
	out_13 <= out_of_13_13;
	out_14 <= out_of_14_13;
	out_15 <= out_of_15_13;
	end
  5'b01111 : 	
	begin
	out_0 <=   out_of_0_12; 
	out_1 <=   out_of_1_12; 
	out_2 <=   out_of_2_12; 
	out_3 <=   out_of_3_12; 
	out_4 <=   out_of_4_12; 
	out_5 <=   out_of_5_12; 
	out_6 <=   out_of_6_12; 
	out_7 <=   out_of_7_12; 
	out_8 <=   out_of_8_12; 
	out_9 <=   out_of_9_12; 
	out_10 <= out_of_10_12;
	out_11 <= out_of_11_12;
	out_12 <= out_of_12_12;
	out_13 <= out_of_13_12;
	out_14 <= out_of_14_12;
	out_15 <= out_of_15_12;
	end




  5'b10000 : 
	begin
	out_0 <=   out_of_0_11; 
	out_1 <=   out_of_1_11; 
	out_2 <=   out_of_2_11; 
	out_3 <=   out_of_3_11; 
	out_4 <=   out_of_4_11; 
	out_5 <=   out_of_5_11; 
	out_6 <=   out_of_6_11; 
	out_7 <=   out_of_7_11; 
	out_8 <=   out_of_8_11; 
	out_9 <=   out_of_9_11; 
	out_10 <= out_of_10_11;
	out_11 <= out_of_11_11;
	out_12 <= out_of_12_11;
	out_13 <= out_of_13_11;
	out_14 <= out_of_14_11;
	out_15 <= out_of_15_11;
	end

  5'b10001 : 	
	begin
	out_0 <=   out_of_0_10; 
	out_1 <=   out_of_1_10; 
	out_2 <=   out_of_2_10; 
	out_3 <=   out_of_3_10; 
	out_4 <=   out_of_4_10; 
	out_5 <=   out_of_5_10; 
	out_6 <=   out_of_6_10; 
	out_7 <=   out_of_7_10; 
	out_8 <=   out_of_8_10; 
	out_9 <=   out_of_9_10; 
	out_10 <= out_of_10_10;
	out_11 <= out_of_11_10;
	out_12 <= out_of_12_10;
	out_13 <= out_of_13_10;
	out_14 <= out_of_14_10;
	out_15 <= out_of_15_10;
	end

  5'b10010 : 	
	begin
	out_0 <=   out_of_0_9; 
	out_1 <=   out_of_1_9; 
	out_2 <=   out_of_2_9; 
	out_3 <=   out_of_3_9; 
	out_4 <=   out_of_4_9; 
	out_5 <=   out_of_5_9; 
	out_6 <=   out_of_6_9; 
	out_7 <=   out_of_7_9; 
	out_8 <=   out_of_8_9; 
	out_9 <=   out_of_9_9; 
	out_10 <= out_of_10_9;
	out_11 <= out_of_11_9;
	out_12 <= out_of_12_9;
	out_13 <= out_of_13_9;
	out_14 <= out_of_14_9;
	out_15 <= out_of_15_9;
	end
  5'b10011 : 	
	begin
	out_0 <=   out_of_0_8; 
	out_1 <=   out_of_1_8; 
	out_2 <=   out_of_2_8; 
	out_3 <=   out_of_3_8; 
	out_4 <=   out_of_4_8; 
	out_5 <=   out_of_5_8; 
	out_6 <=   out_of_6_8; 
	out_7 <=   out_of_7_8; 
	out_8 <=   out_of_8_8; 
	out_9 <=   out_of_9_8; 
	out_10 <= out_of_10_8;
	out_11 <= out_of_11_8;
	out_12 <= out_of_12_8;
	out_13 <= out_of_13_8;
	out_14 <= out_of_14_8;
	out_15 <= out_of_15_8;
	end
  5'b10100 : 	
	begin
	out_0 <=   out_of_0_7; 
	out_1 <=   out_of_1_7; 
	out_2 <=   out_of_2_7; 
	out_3 <=   out_of_3_7; 
	out_4 <=   out_of_4_7; 
	out_5 <=   out_of_5_7; 
	out_6 <=   out_of_6_7; 
	out_7 <=   out_of_7_7; 
	out_8 <=   out_of_8_7; 
	out_9 <=   out_of_9_7; 
	out_10 <= out_of_10_7;
	out_11 <= out_of_11_7;
	out_12 <= out_of_12_7;
	out_13 <= out_of_13_7;
	out_14 <= out_of_14_7;
	out_15 <= out_of_15_7;
	end
  5'b10101 : 	
	begin
	out_0 <=   out_of_0_6; 
	out_1 <=   out_of_1_6; 
	out_2 <=   out_of_2_6; 
	out_3 <=   out_of_3_6; 
	out_4 <=   out_of_4_6; 
	out_5 <=   out_of_5_6; 
	out_6 <=   out_of_6_6; 
	out_7 <=   out_of_7_6; 
	out_8 <=   out_of_8_6; 
	out_9 <=   out_of_9_6; 
	out_10 <= out_of_10_6;
	out_11 <= out_of_11_6;
	out_12 <= out_of_12_6;
	out_13 <= out_of_13_6;
	out_14 <= out_of_14_6;
	out_15 <= out_of_15_6;
	end
  5'b10110 : 	
	begin
	out_0 <=   out_of_0_5; 
	out_1 <=   out_of_1_5; 
	out_2 <=   out_of_2_5; 
	out_3 <=   out_of_3_5; 
	out_4 <=   out_of_4_5; 
	out_5 <=   out_of_5_5; 
	out_6 <=   out_of_6_5; 
	out_7 <=   out_of_7_5; 
	out_8 <=   out_of_8_5; 
	out_9 <=   out_of_9_5; 
	out_10 <= out_of_10_5;
	out_11 <= out_of_11_5;
	out_12 <= out_of_12_5;
	out_13 <= out_of_13_5;
	out_14 <= out_of_14_5;
	out_15 <= out_of_15_5;
	end
  5'b10111 : 	
	begin
	out_0 <=   out_of_0_4; 
	out_1 <=   out_of_1_4; 
	out_2 <=   out_of_2_4; 
	out_3 <=   out_of_3_4; 
	out_4 <=   out_of_4_4; 
	out_5 <=   out_of_5_4; 
	out_6 <=   out_of_6_4; 
	out_7 <=   out_of_7_4; 
	out_8 <=   out_of_8_4; 
	out_9 <=   out_of_9_4; 
	out_10 <= out_of_10_4;
	out_11 <= out_of_11_4;
	out_12 <= out_of_12_4;
	out_13 <= out_of_13_4;
	out_14 <= out_of_14_4;
	out_15 <= out_of_15_4;
	end


5'b11000 : 
	begin
	out_0 <=   out_of_0_3; 
	out_1 <=   out_of_1_3; 
	out_2 <=   out_of_2_3; 
	out_3 <=   out_of_3_3; 
	out_4 <=   out_of_4_3; 
	out_5 <=   out_of_5_3; 
	out_6 <=   out_of_6_3; 
	out_7 <=   out_of_7_3; 
	out_8 <=   out_of_8_3; 
	out_9 <=   out_of_9_3; 
	out_10 <= out_of_10_3;
	out_11 <= out_of_11_3;
	out_12 <= out_of_12_3;
	out_13 <= out_of_13_3;
	out_14 <= out_of_14_3;
	out_15 <= out_of_15_3;
	end

  5'b11001 : 	
	begin
	out_0 <=   out_of_0_2; 
	out_1 <=   out_of_1_2; 
	out_2 <=   out_of_2_2; 
	out_3 <=   out_of_3_2; 
	out_4 <=   out_of_4_2; 
	out_5 <=   out_of_5_2; 
	out_6 <=   out_of_6_2; 
	out_7 <=   out_of_7_2; 
	out_8 <=   out_of_8_2; 
	out_9 <=   out_of_9_2; 
	out_10 <= out_of_10_2;
	out_11 <= out_of_11_2;
	out_12 <= out_of_12_2;
	out_13 <= out_of_13_2;
	out_14 <= out_of_14_2;
	out_15 <= out_of_15_2;
	end

  5'b11010 : 	
	begin
	out_0 <=   out_of_0_1; 
	out_1 <=   out_of_1_1; 
	out_2 <=   out_of_2_1; 
	out_3 <=   out_of_3_1; 
	out_4 <=   out_of_4_1; 
	out_5 <=   out_of_5_1; 
	out_6 <=   out_of_6_1; 
	out_7 <=   out_of_7_1; 
	out_8 <=   out_of_8_1; 
	out_9 <=   out_of_9_1; 
	out_10 <= out_of_10_1;
	out_11 <= out_of_11_1;
	out_12 <= out_of_12_1;
	out_13 <= out_of_13_1;
	out_14 <= out_of_14_1;
	out_15 <= out_of_15_1;
	end
  5'b11011 : 	
	begin
	out_0 <=   out_of_0_0; 
	out_1 <=   out_of_1_0; 
	out_2 <=   out_of_2_0; 
	out_3 <=   out_of_3_0; 
	out_4 <=   out_of_4_0; 
	out_5 <=   out_of_5_0; 
	out_6 <=   out_of_6_0; 
	out_7 <=   out_of_7_0; 
	out_8 <=   out_of_8_0; 
	out_9 <=   out_of_9_0; 
	out_10 <= out_of_10_0;
	out_11 <= out_of_11_0;
	out_12 <= out_of_12_0;
	out_13 <= out_of_13_0;
	out_14 <= out_of_14_0;
	out_15 <= out_of_15_0;
	end
  default : begin
	out_0 <=  0; 
	out_1 <=  0; 
	out_2 <=  0; 
	out_3 <=  0; 
	out_4 <=  0; 
	out_5 <=  0; 
	out_6 <=  0; 
	out_7 <=  0; 
	out_8 <=  0; 
	out_9 <=  0; 
	out_10 <= 0;
	out_11 <= 0;
	out_12 <= 0;
	out_13 <= 0;
	out_14 <= 0;
	out_15 <= 0;
	end
endcase

endmodule